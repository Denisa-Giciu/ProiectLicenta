--componenta deplasator la stanga(shift left)
--este folosita pentru deplasarile la stanga ale bitilor

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity shifter is
	generic (n1: natural:= 32; n2: natural:= 32; k: natural:= 2);
	port (
		x: in std_logic_vector(n1-1 downto 0);
		y: out std_logic_vector(n2-1 downto 0)
	);
end entity;

architecture beh of shifter is
	signal temp: std_logic_vector(n2-1 downto 0);

	begin
	temp <= std_logic_vector(resize(unsigned(x), n2)); --este necesar in cazul maririi sau a micsorarii numarului de biti
	y <= std_logic_vector(shift_left(signed(temp), k));
end beh;